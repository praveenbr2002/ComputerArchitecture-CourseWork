
module tb();

reg [63:0] A,B;
wire [63:0] Product;
wire Cout;

DPFPM F1 (A,B,Product);

initial
begin
    A=64'b0100000010010011010010100100010101101101010111001111101010101101; // 1234.5678
	B=64'b0100000010110110001011100001111110010111001001000111010001010100; // 5678.1234
	#10
	
	
    A=64'b0100000010010011010010100100010101101101010111001111101010101101; // 1234.5678
	B=64'b0; // Zero
	#10
	
    A=64'b01111_1111_1110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_000; // infinity
	B=64'b1100000010110110001011100001111110010111001001000111010001010100; // 5678.1234
	#10
	
	$finish;
end

initial
begin
  $monitor(" %b * %b \n= %b\n", A,B,Product);
end

endmodule
